import bitutils::*;
import bundle::*;
import micro_ops::*;
import csr_def::*;
import exception::*;
