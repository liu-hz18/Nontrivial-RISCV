// I-TLB
import bitutils::*;
import bundle::*;
import csr_def::*;
