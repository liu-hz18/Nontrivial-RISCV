import bitutils::*;
import bundle::*;

module BusSRAM (
    input clk, rst

    // 
);

endmodule

