// 3-pipelined inst-cache
import bitutils::*;
import bundle::*;

module ICache #(
    parameter NAME = "ICACHE"

) (
    input clk, rst,

    input logic flush


);



endmodule
