import bitutils::*;
import bundle::*;
