import bitutils::*;
